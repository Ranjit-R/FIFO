// package fifo_pkg;
//   import uvm_pkg::*;
//   `include "uvm_macros.svh"

//   // Sequence items and sequences
// //   `include "fifo_write_sequence_item.sv"
// //   `include "fifo_read_sequence_item.sv"
//   `include "fifo_sequence_item.sv"
//   `include "fifo_sequence.sv"

//   // Sequencers
//   `include "fifo_sequencer.sv"

//   // Drivers
//   `include "fifo_write_driver.sv"
//   `include "fifo_read_driver.sv"

//   // Monitors
//   `include "fifo_write_monitor.sv"
//   `include "fifo_read_monitor.sv"

//   // Agents
//   `include "fifo_write_agent.sv"
//   `include "fifo_read_agent.sv"

//   // Scoreboard
//   `include "fifo_scoreboard.sv"

//   // (Optional) Functional Coverage
//   // `include "fifo_func_cov.sv"

//   // Environment and Test
//   `include "fifo_env.sv"
//   `include "fifo_test.sv"

// endpackage

