`define ADDR_WIDTH 4
`define DATA_WIDTH 8

`define no_trans 10000 


